library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use model.explicit_params.ALL;
package model_structure is
    constant CONFIG_WIDTH : integer := 168;
    constant AB_PARAMS : T_MODEL_PARAMS := (10, 16, 1, CONFIG_WIDTH);

    subtype T_CONFIGURATION is std_logic_vector(CONFIG_WIDTH-1 downto 0);
    pure function config2lv(c : T_CONFIGURATION) return std_logic_vector;
    pure function lv2config(lv : std_logic_vector) return T_CONFIGURATION;
end package;

package body model_structure is
    pure function config2lv(c : T_CONFIGURATION) return std_logic_vector is
    begin
    	return std_logic_vector(c);
    end function;

    pure function lv2config(lv : std_logic_vector) return T_CONFIGURATION is
    begin
        return T_CONFIGURATION(lv);
    end function;
end package body;

-- /Users/ciprian/Playfield/repositories/plugTEAM/plug-editor-fx/exemples/AliceBobMeetPeterson.fcr state-space
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.explicit_structure.ALL;
use WORK.model_structure.ALL;
package model is
	constant AB_MODEL : T_EXPLICIT := (
		states => (
			0 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000001_00000000_00000000",
			1 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000",
			2 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000001_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000",
			3 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000",
			4 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000",
			5 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000001_00000000_00000011_00000000_00000000",
			6 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000001_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000",
			7 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000001_00000001_00000000_00000000_00000000_00000010_00000000_00000011_00000000_00000000",
			8 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000001_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000",
			9 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000001_00000000_00000000"		),
		initial => (0 => 0),
		fanout => (
			3, 1			-- fanout(0)
			, 2, 5			-- fanout(1)
			, 7			-- fanout(2)
			, 4, 8			-- fanout(3)
			, 9, 6			-- fanout(4)
			, 7, 0			-- fanout(5)
			, 1			-- fanout(6)
			, 3			-- fanout(7)
			, 6			-- fanout(8)
			, 3, 1			-- fanout(9)
		),
		fanout_base => (0, 2, 4, 5, 7, 9, 11, 12, 13, 14, 16)
);
end package;
