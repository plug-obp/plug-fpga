-- /Users/ciprian/Playfield/repositories/beem-benchmark/fiacre-version/bakery/generated_files/bakery_1.fcr state-space
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use WORK.explicit_structure.ALL;
use WORK.model_structure.ALL;
package model is
	constant AB_MODEL : T_EXPLICIT := (
		states => (
			0 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			2 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			3 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			4 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			5 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			6 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			7 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			8 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			9 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			10 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			11 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			12 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			13 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			14 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			15 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			16 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			17 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			18 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			19 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			20 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			21 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			22 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			23 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			24 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			25 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			26 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			27 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			28 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			29 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			30 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			31 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			32 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			33 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			34 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			35 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			36 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			37 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			38 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			39 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			40 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			41 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			42 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			43 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			44 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			45 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			46 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			47 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			48 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			49 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			50 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			51 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			52 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			53 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			54 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			55 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			56 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			57 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			58 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			59 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			60 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			61 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			62 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			63 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			64 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			65 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			66 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			67 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			68 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			69 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			70 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			71 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			72 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			73 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			74 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			75 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			76 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			77 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			78 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			79 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			80 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			81 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			82 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			83 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			84 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			85 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			86 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			87 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			88 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			89 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			90 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			91 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			92 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			93 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			94 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			95 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			96 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			97 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			98 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			99 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			100 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			101 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			102 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			103 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			104 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			105 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			106 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			107 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			108 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			109 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			110 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			111 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			112 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			113 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			114 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			115 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			116 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			117 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			118 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			119 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			120 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			121 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			122 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			123 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			124 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			125 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			126 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			127 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			128 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			129 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			130 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			131 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			132 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			133 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			134 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			135 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			136 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			137 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			138 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			139 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			140 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			141 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			142 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			143 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			144 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			145 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			146 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			147 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			148 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			149 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			150 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			151 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			152 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			153 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			154 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			155 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			156 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			157 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			158 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			159 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			160 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			161 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			162 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			163 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			164 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			165 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			166 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			167 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			168 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			169 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			170 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			171 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			172 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			173 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			174 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			175 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			176 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			177 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			178 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			179 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			180 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			181 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			182 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			183 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			184 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			185 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			186 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			187 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			188 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			189 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			190 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			191 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			192 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			193 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			194 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			195 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			196 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			197 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			198 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			199 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			200 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			201 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			202 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			203 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			204 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			205 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			206 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			207 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			208 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			209 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			210 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			211 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			212 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			213 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			214 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			215 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			216 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			217 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			218 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			219 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			220 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			221 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			222 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			223 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			224 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			225 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			226 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			227 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			228 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			229 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			230 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			231 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			232 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			233 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			234 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			235 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			236 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			237 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			238 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			239 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			240 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			241 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			242 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			243 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			244 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			245 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			246 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			247 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			248 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			249 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			250 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			251 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			252 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			253 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			254 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			255 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			256 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			257 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			258 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			259 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			260 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			261 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			262 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			263 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			264 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			265 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			266 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			267 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			268 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			269 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			270 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			271 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			272 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			273 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			274 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			275 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			276 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			277 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			278 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			279 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			280 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			281 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			282 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			283 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			284 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			285 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			286 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			287 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			288 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			289 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			290 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			291 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			292 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			293 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			294 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			295 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			296 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			297 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			298 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			299 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			300 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			301 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			302 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			303 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			304 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			305 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			306 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			307 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			308 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			309 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			310 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			311 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			312 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			313 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			314 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			315 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			316 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			317 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			318 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			319 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			320 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			321 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			322 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			323 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			324 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			325 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			326 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			327 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			328 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			329 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			330 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			331 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			332 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			333 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			334 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			335 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			336 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			337 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			338 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			339 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			340 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			341 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			342 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			343 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			344 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			345 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			346 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			347 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			348 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			349 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			350 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			351 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			352 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			353 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			354 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			355 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			356 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			357 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			358 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			359 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			360 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			361 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			362 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			363 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			364 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			365 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			366 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			367 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			368 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			369 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			370 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			371 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			372 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			373 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			374 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			375 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			376 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			377 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			378 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			379 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			380 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			381 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			382 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			383 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			384 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			385 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			386 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			387 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			388 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			389 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			390 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			391 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			392 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			393 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			394 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			395 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			396 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			397 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			398 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			399 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			400 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			401 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			402 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			403 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			404 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			405 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			406 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			407 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			408 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			409 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			410 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			411 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			412 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			413 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			414 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			415 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			416 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			417 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			418 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			419 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			420 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			421 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			422 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			423 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			424 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			425 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			426 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			427 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			428 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			429 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			430 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			431 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			432 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			433 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			434 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			435 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			436 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			437 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			438 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			439 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			440 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			441 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			442 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			443 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			444 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			445 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			446 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			447 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			448 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			449 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			450 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			451 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			452 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			453 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			454 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			455 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			456 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			457 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			458 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			459 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			460 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			461 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			462 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			463 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			464 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			465 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			466 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			467 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			468 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			469 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			470 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			471 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			472 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			473 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			474 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			475 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			476 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			477 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			478 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			479 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			480 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			481 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			482 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			483 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			484 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			485 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			486 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			487 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			488 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			489 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			490 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			491 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			492 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			493 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			494 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			495 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			496 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			497 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			498 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			499 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			500 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			501 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			502 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			503 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			504 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			505 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			506 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			507 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			508 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			509 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			510 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			511 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			512 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			513 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			514 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			515 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			516 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			517 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			518 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			519 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			520 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			521 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			522 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			523 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			524 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			525 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			526 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			527 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			528 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			529 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			530 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			531 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			532 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			533 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			534 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			535 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			536 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			537 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			538 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			539 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			540 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			541 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			542 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			543 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			544 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			545 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			546 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			547 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			548 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			549 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			550 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			551 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			552 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			553 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			554 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			555 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			556 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			557 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			558 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			559 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			560 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			561 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			562 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			563 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			564 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			565 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			566 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			567 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			568 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			569 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			570 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			571 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			572 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			573 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			574 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			575 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			576 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			577 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			578 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			579 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			580 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			581 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			582 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			583 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			584 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			585 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			586 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			587 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			588 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			589 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			590 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			591 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			592 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			593 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			594 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			595 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			596 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			597 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			598 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			599 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			600 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			601 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			602 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			603 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			604 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			605 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			606 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			607 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			608 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			609 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			610 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			611 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			612 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			613 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			614 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			615 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			616 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			617 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			618 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			619 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			620 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			621 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			622 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			623 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			624 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			625 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			626 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			627 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			628 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			629 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			630 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			631 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			632 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			633 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			634 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			635 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			636 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			637 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			638 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			639 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			640 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			641 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			642 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			643 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			644 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			645 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			646 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			647 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			648 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			649 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			650 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			651 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			652 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			653 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			654 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			655 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			656 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			657 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			658 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			659 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			660 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			661 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			662 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			663 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			664 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			665 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			666 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			667 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			668 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			669 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			670 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			671 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			672 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			673 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			674 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			675 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			676 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			677 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			678 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			679 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			680 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			681 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			682 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			683 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			684 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			685 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			686 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			687 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			688 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			689 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			690 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			691 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			692 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			693 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			694 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			695 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			696 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			697 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			698 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			699 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			700 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			701 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			702 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			703 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			704 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			705 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			706 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			707 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			708 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			709 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			710 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			711 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			712 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			713 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			714 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			715 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			716 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			717 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			718 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			719 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			720 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			721 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			722 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			723 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			724 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			725 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			726 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			727 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			728 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			729 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			730 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			731 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			732 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			733 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			734 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			735 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			736 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			737 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			738 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			739 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			740 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			741 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			742 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			743 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			744 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			745 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			746 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			747 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			748 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			749 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			750 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			751 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			752 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			753 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			754 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			755 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			756 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			757 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			758 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			759 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			760 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			761 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			762 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			763 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			764 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			765 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			766 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			767 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			768 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			769 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			770 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			771 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			772 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			773 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			774 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			775 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			776 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			777 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			778 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			779 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			780 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			781 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			782 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			783 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			784 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			785 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			786 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			787 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			788 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			789 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			790 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			791 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			792 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			793 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			794 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			795 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			796 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			797 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			798 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			799 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			800 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			801 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			802 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			803 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			804 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			805 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			806 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			807 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			808 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			809 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			810 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			811 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			812 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			813 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			814 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			815 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			816 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			817 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			818 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			819 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			820 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			821 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			822 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			823 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			824 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			825 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			826 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			827 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			828 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			829 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			830 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			831 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			832 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			833 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			834 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			835 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			836 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			837 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			838 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			839 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			840 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			841 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			842 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			843 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			844 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			845 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			846 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			847 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			848 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			849 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			850 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			851 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			852 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			853 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			854 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			855 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			856 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			857 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			858 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			859 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			860 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			861 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			862 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			863 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			864 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			865 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			866 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			867 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			868 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			869 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			870 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			871 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			872 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			873 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			874 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			875 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			876 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			877 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			878 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			879 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			880 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			881 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			882 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			883 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			884 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			885 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			886 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			887 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			888 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			889 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			890 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			891 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			892 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			893 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			894 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			895 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			896 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			897 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			898 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			899 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			900 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			901 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			902 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			903 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			904 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			905 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			906 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			907 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			908 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			909 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			910 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			911 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			912 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			913 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			914 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			915 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			916 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			917 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			918 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			919 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			920 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			921 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			922 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			923 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			924 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			925 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			926 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			927 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			928 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			929 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			930 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			931 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			932 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			933 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			934 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			935 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			936 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			937 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			938 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			939 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			940 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			941 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			942 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			943 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			944 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			945 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			946 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			947 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			948 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			949 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			950 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			951 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			952 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			953 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			954 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			955 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			956 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			957 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			958 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			959 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			960 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			961 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			962 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			963 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			964 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			965 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			966 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			967 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			968 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			969 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			970 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			971 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			972 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			973 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			974 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			975 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			976 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			977 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			978 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			979 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			980 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			981 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			982 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			983 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			984 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			985 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			986 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			987 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			988 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			989 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			990 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			991 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			992 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			993 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			994 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			995 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			996 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			997 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			998 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			999 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1000 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1001 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1002 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1003 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1004 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1005 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1006 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1007 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1008 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1009 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1010 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1011 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1012 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1013 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1014 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1015 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1016 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1017 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1018 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1019 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1020 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1021 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1022 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1023 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1024 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1025 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1026 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1027 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1028 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1029 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1030 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1031 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1032 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1033 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1034 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1035 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1036 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1037 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1038 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1039 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1040 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1041 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1042 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1043 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1044 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1045 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1046 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1047 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1048 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1049 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1050 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1051 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1052 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1053 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1054 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1055 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1056 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1057 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1058 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1059 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1060 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1061 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1062 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1063 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1064 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1065 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1066 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1067 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1068 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1069 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1070 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1071 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1072 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1073 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1074 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1075 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1076 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1077 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1078 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1079 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1080 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1081 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1082 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1083 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1084 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1085 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1086 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1087 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1088 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1089 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1090 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1091 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1092 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1093 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1094 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1095 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1096 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1097 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1098 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1099 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1100 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1101 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1102 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1103 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1104 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1105 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1106 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1107 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1108 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1109 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1110 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1111 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1112 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1113 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1114 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1115 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1116 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1117 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1118 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1119 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1120 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1121 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1122 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1123 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1124 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1125 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1126 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1127 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1128 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1129 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1130 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1131 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1132 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1133 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1134 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1135 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1136 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1137 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1138 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1139 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1140 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1141 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1142 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1143 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1144 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1145 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1146 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1147 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1148 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1149 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1150 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1151 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1152 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1153 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1154 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1155 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1156 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1157 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1158 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1159 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1160 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1161 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1162 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1163 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1164 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1165 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1166 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1167 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1168 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1169 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1170 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1171 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1172 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1173 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1174 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1175 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1176 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1177 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1178 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1179 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1180 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1181 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1182 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1183 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1184 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1185 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1186 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1187 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1188 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1189 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1190 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1191 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1192 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1193 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1194 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1195 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1196 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1197 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1198 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1199 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1200 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1201 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1202 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1203 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1204 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1205 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1206 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1207 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1208 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1209 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1210 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1211 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1212 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1213 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1214 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1215 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1216 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1217 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1218 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1219 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1220 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1221 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1222 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1223 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1224 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1225 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1226 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1227 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1228 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1229 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1230 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1231 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1232 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1233 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1234 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1235 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1236 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1237 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1238 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1239 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1240 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1241 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1242 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1243 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1244 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1245 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1246 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1247 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1248 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1249 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1250 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1251 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1252 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1253 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1254 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1255 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1256 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1257 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1258 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1259 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1260 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1261 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1262 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1263 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1264 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1265 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1266 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1267 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1268 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1269 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1270 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1271 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1272 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1273 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1274 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1275 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1276 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1277 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1278 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1279 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1280 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1281 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1282 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1283 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1284 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1285 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1286 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1287 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1288 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1289 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1290 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1291 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1292 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1293 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1294 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1295 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1296 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1297 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1298 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1299 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1300 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1301 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1302 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1303 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1304 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1305 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1306 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1307 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1308 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1309 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1310 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1311 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1312 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1313 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1314 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1315 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1316 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1317 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1318 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1319 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1320 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1321 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1322 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1323 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1324 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1325 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1326 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1327 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1328 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1329 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1330 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1331 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1332 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1333 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1334 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1335 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1336 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1337 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1338 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1339 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1340 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1341 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1342 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1343 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1344 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1345 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1346 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1347 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1348 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1349 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1350 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1351 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1352 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1353 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1354 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1355 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1356 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1357 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1358 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1359 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1360 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1361 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1362 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1363 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1364 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1365 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1366 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1367 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1368 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1369 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1370 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1371 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1372 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1373 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1374 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1375 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1376 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1377 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1378 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1379 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1380 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1381 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1382 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1383 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1384 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1385 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1386 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1387 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1388 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1389 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1390 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1391 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1392 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1393 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1394 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1395 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1396 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1397 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1398 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1399 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1400 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1401 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1402 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1403 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1404 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1405 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1406 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1407 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1408 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1409 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1410 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1411 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1412 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1413 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1414 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1415 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1416 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1417 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1418 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1419 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1420 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1421 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1422 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1423 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1424 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1425 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1426 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1427 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1428 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1429 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1430 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1431 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1432 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1433 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1434 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1435 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000",
			1436 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1437 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1438 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1439 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1440 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1441 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1442 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1443 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1444 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1445 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1446 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1447 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1448 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1449 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1450 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1451 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1452 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1453 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1454 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1455 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1456 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1457 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1458 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1459 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1460 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1461 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1462 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1463 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1464 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1465 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1466 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1467 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1468 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1469 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1470 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1471 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1472 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1473 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1474 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1475 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1476 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1477 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1478 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1479 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1480 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1481 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1482 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1483 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1484 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1485 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1486 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1487 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000000",
			1488 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000",
			1489 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1490 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1491 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1492 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000010_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000000",
			1493 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1494 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1495 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1496 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000001_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1497 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00001000_00000000_00000000_00000000_00000010_00000000_00000001_00000000_00000000_00000000_00001001_00000000_00000000_00000000_00000000",
			1498 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1499 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000000",
			1500 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000",
			1501 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000110_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000000_00000000_00000101_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000",
			1502 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000100_00000000_00000001_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000011_00000000_00000010_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000",
			1503 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1504 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010_00000000_00000010_00000000_00000000_00000000_00000111_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000",
			1505 => B"00000001_00000011_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001_00000010_00000000_00000000_00000000_00000011_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000011_00000000_00000001_00000000_00000000_00000000_00000010_00000000_00000000_00000000_00000100_00000000_00000000_00000000_00000000_00000000_00000001_00000000_00000000_00000000_00000000"		),
		initial => (0 => 131),
		fanout => (
			1330, 17			-- fanout(0)
			, 286			-- fanout(1)
			, 1069, 287			-- fanout(2)
			, 759, 18			-- fanout(3)
			, 761, 10			-- fanout(4)
			, 14			-- fanout(5)
			, 702, 9			-- fanout(6)
			, 788, 11			-- fanout(7)
			, 37, 326			-- fanout(8)
			, 1113, 285			-- fanout(9)
			, 769, 289			-- fanout(10)
			, 770, 631			-- fanout(11)
			, 96, 266			-- fanout(12)
			, 1320, 315			-- fanout(13)
			, 291			-- fanout(14)
			, 771, 1308			-- fanout(15)
			, 1103, 312			-- fanout(16)
			, 1325			-- fanout(17)
			, 752, 296			-- fanout(18)
			, 1354, 30			-- fanout(19)
			, 425, 938			-- fanout(20)
			, 51, 929			-- fanout(21)
			, 805, 923			-- fanout(22)
			, 358, 29			-- fanout(23)
			, 710, 27			-- fanout(24)
			, 1364, 901			-- fanout(25)
			, 1368, 901			-- fanout(26)
			, 706, 308			-- fanout(27)
			, 407, 938			-- fanout(28)
			, 343, 57			-- fanout(29)
			, 1351, 304			-- fanout(30)
			, 776, 923			-- fanout(31)
			, 328			-- fanout(32)
			, 801			-- fanout(33)
			, 799, 732			-- fanout(34)
			, 938, 303			-- fanout(35)
			, 803, 319			-- fanout(36)
			, 832, 39			-- fanout(37)
			, 122, 299			-- fanout(38)
			, 814, 51			-- fanout(39)
			, 1374, 512			-- fanout(40)
			, 798, 674			-- fanout(41)
			, 301			-- fanout(42)
			, 1310			-- fanout(43)
			, 777, 6			-- fanout(44)
			, 1405, 13			-- fanout(45)
			, 1401			-- fanout(46)
			, 5			-- fanout(47)
			, 1429, 45			-- fanout(48)
			, 772, 64			-- fanout(49)
			, 1430, 46			-- fanout(50)
			, 856, 981			-- fanout(51)
			, 644			-- fanout(52)
			, 105, 8			-- fanout(53)
			, 415, 980			-- fanout(54)
			, 840, 36			-- fanout(55)
			, 648, 190			-- fanout(56)
			, 404, 980			-- fanout(57)
			, 842, 1440			-- fanout(58)
			, 533, 317			-- fanout(59)
			, 830, 33			-- fanout(60)
			, 452, 995			-- fanout(61)
			, 829, 41			-- fanout(62)
			, 647, 772			-- fanout(63)
			, 762, 16			-- fanout(64)
			, 658, 200			-- fanout(65)
			, 150, 53			-- fanout(66)
			, 650, 1459			-- fanout(67)
			, 1394, 323			-- fanout(68)
			, 663, 789			-- fanout(69)
			, 685			-- fanout(70)
			, 1396			-- fanout(71)
			, 800, 84			-- fanout(72)
			, 884			-- fanout(73)
			, 662, 1472			-- fanout(74)
			, 671, 800			-- fanout(75)
			, 665, 216			-- fanout(76)
			, 435, 23			-- fanout(77)
			, 882, 82			-- fanout(78)
			, 675, 1482			-- fanout(79)
			, 844, 97			-- fanout(80)
			, 1449, 1020			-- fanout(81)
			, 850			-- fanout(82)
			, 1480			-- fanout(83)
			, 791, 24			-- fanout(84)
			, 1362, 88			-- fanout(85)
			, 322			-- fanout(86)
			, 858, 7			-- fanout(87)
			, 1332			-- fanout(88)
			, 1303, 43			-- fanout(89)
			, 789, 44			-- fanout(90)
			, 47			-- fanout(91)
			, 854, 981			-- fanout(92)
			, 70			-- fanout(93)
			, 425, 980			-- fanout(94)
			, 1419, 1494			-- fanout(95)
			, 751, 2			-- fanout(96)
			, 862			-- fanout(97)
			, 847, 87			-- fanout(98)
			, 873, 113			-- fanout(99)
			, 536			-- fanout(100)
			, 357			-- fanout(101)
			, 407, 1093			-- fanout(102)
			, 1063			-- fanout(103)
			, 1390, 107			-- fanout(104)
			, 532, 37			-- fanout(105)
			, 877, 110			-- fanout(106)
			, 1384			-- fanout(107)
			, 1474, 235			-- fanout(108)
			, 1476, 40			-- fanout(109)
			, 886			-- fanout(110)
			, 1349, 116			-- fanout(111)
			, 1059, 1047			-- fanout(112)
			, 868			-- fanout(113)
			, 1455, 1020			-- fanout(114)
			, 881, 1500			-- fanout(115)
			, 1365			-- fanout(116)
			, 446, 77			-- fanout(117)
			, 870, 1138			-- fanout(118)
			, 890, 73			-- fanout(119)
			, 529, 58			-- fanout(120)
			, 530, 136			-- fanout(121)
			, 626, 59			-- fanout(122)
			, 839, 1060			-- fanout(123)
			, 346, 415			-- fanout(124)
			, 821, 1055			-- fanout(125)
			, 567, 146			-- fanout(126)
			, 1411, 1111			-- fanout(127)
			, 1077, 112			-- fanout(128)
			, 1497, 71			-- fanout(129)
			, 42			-- fanout(130)
			, 236, 1316			-- fanout(131)
			, 547, 62			-- fanout(132)
			, 538			-- fanout(133)
			, 425, 1093			-- fanout(134)
			, 535, 34			-- fanout(135)
			, 548, 55			-- fanout(136)
			, 766, 1162			-- fanout(137)
			, 522, 132			-- fanout(138)
			, 369, 124			-- fanout(139)
			, 361, 418			-- fanout(140)
			, 409, 1093			-- fanout(141)
			, 103			-- fanout(142)
			, 372, 52			-- fanout(143)
			, 628, 1068			-- fanout(144)
			, 1465, 1164			-- fanout(145)
			, 544, 405			-- fanout(146)
			, 101			-- fanout(147)
			, 1367, 66			-- fanout(148)
			, 540, 100			-- fanout(149)
			, 542, 105			-- fanout(150)
			, 524, 133			-- fanout(151)
			, 178			-- fanout(152)
			, 1489			-- fanout(153)
			, 843, 125			-- fanout(154)
			, 371, 56			-- fanout(155)
			, 1357			-- fanout(156)
			, 378, 67			-- fanout(157)
			, 373, 63			-- fanout(158)
			, 588, 1079			-- fanout(159)
			, 384, 65			-- fanout(160)
			, 1136, 95			-- fanout(161)
			, 1135, 882			-- fanout(162)
			, 1137, 274			-- fanout(163)
			, 390, 140			-- fanout(164)
			, 590, 180			-- fanout(165)
			, 380, 425			-- fanout(166)
			, 381, 69			-- fanout(167)
			, 392, 76			-- fanout(168)
			, 387, 74			-- fanout(169)
			, 394, 75			-- fanout(170)
			, 1226, 704			-- fanout(171)
			, 1505, 48			-- fanout(172)
			, 638, 144			-- fanout(173)
			, 563, 1308			-- fanout(174)
			, 83			-- fanout(175)
			, 1484, 68			-- fanout(176)
			, 393, 79			-- fanout(177)
			, 93			-- fanout(178)
			, 1229, 704			-- fanout(179)
			, 555, 98			-- fanout(180)
			, 1486, 410			-- fanout(181)
			, 1273, 704			-- fanout(182)
			, 1483, 172			-- fanout(183)
			, 1270, 704			-- fanout(184)
			, 1398, 1111			-- fanout(185)
			, 1490, 1078			-- fanout(186)
			, 287, 641			-- fanout(187)
						-- fanout(188)
			, 690, 228			-- fanout(189)
			, 760			-- fanout(190)
			, 1185			-- fanout(191)
			, 7, 499			-- fanout(192)
			, 768, 460			-- fanout(193)
			, 994, 839			-- fanout(194)
			, 106			-- fanout(195)
			, 501			-- fanout(196)
			, 945, 468			-- fanout(197)
			, 967, 438			-- fanout(198)
			, 339, 189			-- fanout(199)
			, 773			-- fanout(200)
			, 956			-- fanout(201)
			, 1, 440			-- fanout(202)
			, 784, 474			-- fanout(203)
			, 954, 198			-- fanout(204)
			, 702, 219			-- fanout(205)
			, 990, 194			-- fanout(206)
			, 149			-- fanout(207)
			, 727, 479			-- fanout(208)
			, 303, 487			-- fanout(209)
			, 309, 1151			-- fanout(210)
			, 982			-- fanout(211)
			, 988, 489			-- fanout(212)
			, 38, 488			-- fanout(213)
			, 1029, 212			-- fanout(214)
			, 992, 220			-- fanout(215)
			, 790			-- fanout(216)
			, 1032, 211			-- fanout(217)
			, 737			-- fanout(218)
			, 1113, 486			-- fanout(219)
			, 1003, 1128			-- fanout(220)
			, 1010, 456			-- fanout(221)
			, 485			-- fanout(222)
			, 983, 465			-- fanout(223)
			, 222			-- fanout(224)
			, 494			-- fanout(225)
			, 1020, 477			-- fanout(226)
			, 1023, 496			-- fanout(227)
			, 368, 1181			-- fanout(228)
			, 36, 519			-- fanout(229)
			, 470			-- fanout(230)
			, 55, 229			-- fanout(231)
			, 1056, 227			-- fanout(232)
			, 225			-- fanout(233)
			, 62, 239			-- fanout(234)
			, 60, 242			-- fanout(235)
			, 810, 1403			-- fanout(236)
			, 1042, 511			-- fanout(237)
			, 42, 482			-- fanout(238)
			, 41, 854			-- fanout(239)
			, 1013, 237			-- fanout(240)
			, 32, 483			-- fanout(241)
			, 33			-- fanout(242)
			, 1154			-- fanout(243)
			, 254			-- fanout(244)
			, 86, 493			-- fanout(245)
			, 97			-- fanout(246)
			, 1336, 1212			-- fanout(247)
			, 1085, 1203			-- fanout(248)
			, 87, 192			-- fanout(249)
			, 462, 230			-- fanout(250)
			, 317, 1005			-- fanout(251)
			, 1063, 1203			-- fanout(252)
			, 414, 199			-- fanout(253)
			, 196			-- fanout(254)
			, 298			-- fanout(255)
			, 450, 253			-- fanout(256)
			, 73			-- fanout(257)
			, 1008, 273			-- fanout(258)
			, 1011, 1204			-- fanout(259)
			, 119, 257			-- fanout(260)
			, 1078, 221			-- fanout(261)
			, 116			-- fanout(262)
			, 1108			-- fanout(263)
			, 1109, 215			-- fanout(264)
			, 1076, 206			-- fanout(265)
			, 2, 187			-- fanout(266)
			, 98, 249			-- fanout(267)
			, 754, 1234			-- fanout(268)
			, 88			-- fanout(269)
			, 1322, 1212			-- fanout(270)
			, 340			-- fanout(271)
			, 85, 269			-- fanout(272)
			, 989, 1211			-- fanout(273)
			, 80, 246			-- fanout(274)
			, 104, 295			-- fanout(275)
			, 1105, 1248			-- fanout(276)
			, 99, 283			-- fanout(277)
			, 708, 1248			-- fanout(278)
			, 130, 238			-- fanout(279)
			, 132, 234			-- fanout(280)
			, 35, 209			-- fanout(281)
			, 136, 231			-- fanout(282)
			, 113			-- fanout(283)
			, 789, 297			-- fanout(284)
			, 1030, 259			-- fanout(285)
			, 165			-- fanout(286)
			, 1001, 366			-- fanout(287)
			, 1123, 263			-- fanout(288)
			, 1121, 265			-- fanout(289)
			, 1112, 214			-- fanout(290)
			, 255			-- fanout(291)
			, 111, 262			-- fanout(292)
			, 1031, 1236			-- fanout(293)
			, 1094, 290			-- fanout(294)
			, 107			-- fanout(295)
			, 1124, 264			-- fanout(296)
			, 777, 205			-- fanout(297)
			, 127, 1282			-- fanout(298)
			, 59, 251			-- fanout(299)
			, 743, 604			-- fanout(300)
			, 1089			-- fanout(301)
			, 174, 1485			-- fanout(302)
			, 1271, 243			-- fanout(303)
			, 138, 280			-- fanout(304)
			, 714, 232			-- fanout(305)
			, 121, 282			-- fanout(306)
			, 705, 305			-- fanout(307)
			, 1044, 293			-- fanout(308)
			, 1197, 1294			-- fanout(309)
			, 1217, 1302			-- fanout(310)
			, 165, 331			-- fanout(311)
			, 1095, 258			-- fanout(312)
			, 89, 334			-- fanout(313)
			, 725, 1308			-- fanout(314)
			, 159, 1277			-- fanout(315)
			, 765, 1308			-- fanout(316)
			, 838, 1119			-- fanout(317)
			, 764, 1308			-- fanout(318)
			, 726, 300			-- fanout(319)
			, 505, 256			-- fanout(320)
			, 720, 1308			-- fanout(321)
			, 271			-- fanout(322)
			, 1339, 1355			-- fanout(323)
			, 734, 1308			-- fanout(324)
			, 729, 1308			-- fanout(325)
			, 39, 21			-- fanout(326)
			, 185, 1282			-- fanout(327)
			, 1354			-- fanout(328)
			, 724, 1308			-- fanout(329)
			, 425, 1316			-- fanout(330)
			, 180, 267			-- fanout(331)
			, 723, 1308			-- fanout(332)
			, 495			-- fanout(333)
			, 43			-- fanout(334)
			, 1178			-- fanout(335)
			, 1176, 350			-- fanout(336)
			, 1186, 1022			-- fanout(337)
			, 442, 620			-- fanout(338)
			, 1180, 690			-- fanout(339)
			, 1218, 354			-- fanout(340)
			, 1183, 347			-- fanout(341)
			, 408			-- fanout(342)
			, 972, 404			-- fanout(343)
			, 204, 692			-- fanout(344)
			, 747, 638			-- fanout(345)
			, 1386, 1050			-- fanout(346)
			, 1169			-- fanout(347)
			, 1168, 353			-- fanout(348)
			, 1189, 694			-- fanout(349)
			, 1174, 643			-- fanout(350)
			, 619			-- fanout(351)
			, 719, 345			-- fanout(352)
			, 1196			-- fanout(353)
			, 1175			-- fanout(354)
			, 187, 830			-- fanout(355)
			, 436, 687			-- fanout(356)
			, 210, 1363			-- fanout(357)
			, 997, 343			-- fanout(358)
			, 1487			-- fanout(359)
			, 991, 409			-- fanout(360)
			, 1187, 1053			-- fanout(361)
			, 217, 388			-- fanout(362)
			, 214, 382			-- fanout(363)
			, 342			-- fanout(364)
			, 237, 661			-- fanout(365)
			, 1143, 359			-- fanout(366)
			, 1085			-- fanout(367)
			, 1239, 1380			-- fanout(368)
			, 1410, 346			-- fanout(369)
			, 386			-- fanout(370)
			, 1012, 648			-- fanout(371)
			, 1004, 644			-- fanout(372)
			, 1016, 647			-- fanout(373)
			, 1019, 360			-- fanout(374)
			, 469, 38			-- fanout(375)
			, 739, 634			-- fanout(376)
			, 1014, 423			-- fanout(377)
			, 1015, 650			-- fanout(378)
			, 632			-- fanout(379)
			, 948, 1071			-- fanout(380)
			, 1025, 663			-- fanout(381)
			, 212, 670			-- fanout(382)
			, 1200, 337			-- fanout(383)
			, 1018, 658			-- fanout(384)
			, 1224, 335			-- fanout(385)
			, 682			-- fanout(386)
			, 1027, 662			-- fanout(387)
			, 211			-- fanout(388)
			, 209, 637			-- fanout(389)
			, 1201, 361			-- fanout(390)
			, 367			-- fanout(391)
			, 1026, 665			-- fanout(392)
			, 1034, 675			-- fanout(393)
			, 1028, 671			-- fanout(394)
			, 699			-- fanout(395)
			, 1039, 377			-- fanout(396)
			, 251, 1183			-- fanout(397)
			, 980, 651			-- fanout(398)
			, 1264, 1116			-- fanout(399)
			, 252, 1414			-- fanout(400)
			, 240, 365			-- fanout(401)
			, 969, 380			-- fanout(402)
			, 1103, 406			-- fanout(403)
			, 1049, 1403			-- fanout(404)
			, 1228, 1380			-- fanout(405)
			, 1095, 645			-- fanout(406)
			, 1047, 1403			-- fanout(407)
			, 1402			-- fanout(408)
			, 1052, 1403			-- fanout(409)
			, 248, 1414			-- fanout(410)
			, 951			-- fanout(411)
			, 1258			-- fanout(412)
			, 1259, 307			-- fanout(413)
			, 1260, 339			-- fanout(414)
			, 1050, 1403			-- fanout(415)
			, 1055, 1403			-- fanout(416)
			, 1249, 399			-- fanout(417)
			, 1053, 1403			-- fanout(418)
			, 942, 411			-- fanout(419)
			, 708			-- fanout(420)
			, 1068, 1403			-- fanout(421)
			, 1292, 336			-- fanout(422)
			, 1061, 1403			-- fanout(423)
			, 266, 355			-- fanout(424)
			, 1071, 1403			-- fanout(425)
			, 693			-- fanout(426)
			, 1269, 288			-- fanout(427)
			, 911			-- fanout(428)
			, 899, 428			-- fanout(429)
			, 1105			-- fanout(430)
			, 804, 352			-- fanout(431)
			, 420			-- fanout(432)
			, 1283, 1434			-- fanout(433)
			, 1279, 383			-- fanout(434)
			, 1088, 358			-- fanout(435)
			, 976, 455			-- fanout(436)
			, 351			-- fanout(437)
			, 1311, 434			-- fanout(438)
			, 290, 363			-- fanout(439)
			, 286, 311			-- fanout(440)
			, 364			-- fanout(441)
			, 836, 376			-- fanout(442)
			, 828			-- fanout(443)
			, 1477, 369			-- fanout(444)
			, 1296, 422			-- fanout(445)
			, 1096, 435			-- fanout(446)
			, 271, 524			-- fanout(447)
			, 430			-- fanout(448)
			, 1290, 412			-- fanout(449)
			, 1299, 414			-- fanout(450)
			, 441			-- fanout(451)
			, 1277, 1434			-- fanout(452)
			, 1102, 374			-- fanout(453)
			, 1481, 444			-- fanout(454)
			, 940			-- fanout(455)
			, 1307, 585			-- fanout(456)
			, 278, 1462			-- fanout(457)
			, 1280, 390			-- fanout(458)
			, 1011, 1461			-- fanout(459)
			, 1115, 453			-- fanout(460)
			, 391			-- fanout(461)
			, 772, 470			-- fanout(462)
			, 281, 389			-- fanout(463)
			, 1128, 1454			-- fanout(464)
			, 912, 4			-- fanout(465)
			, 1122, 396			-- fanout(466)
			, 1306, 1449			-- fanout(467)
			, 1287, 458			-- fanout(468)
			, 999, 122			-- fanout(469)
			, 762, 403			-- fanout(470)
			, 704, 393			-- fanout(471)
			, 1066, 402			-- fanout(472)
			, 294, 439			-- fanout(473)
			, 707, 466			-- fanout(474)
			, 276, 1462			-- fanout(475)
			, 395			-- fanout(476)
			, 902, 427			-- fanout(477)
			, 250, 490			-- fanout(478)
			, 1075, 472			-- fanout(479)
			, 909, 417			-- fanout(480)
			, 300, 776			-- fanout(481)
			, 301, 1290			-- fanout(482)
			, 328, 19			-- fanout(483)
			, 944, 758			-- fanout(484)
			, 461			-- fanout(485)
			, 1030, 459			-- fanout(486)
			, 243			-- fanout(487)
			, 299, 397			-- fanout(488)
			, 900, 467			-- fanout(489)
			, 230			-- fanout(490)
			, 318, 1485			-- fanout(491)
			, 316, 1485			-- fanout(492)
			, 322, 447			-- fanout(493)
			, 503			-- fanout(494)
			, 930, 505			-- fanout(495)
			, 931, 484			-- fanout(496)
			, 314, 1485			-- fanout(497)
			, 12, 424			-- fanout(498)
			, 11, 805			-- fanout(499)
			, 15, 1485			-- fanout(500)
			, 432			-- fanout(501)
			, 270, 1484			-- fanout(502)
			, 448			-- fanout(503)
			, 949, 413			-- fanout(504)
			, 950, 450			-- fanout(505)
			, 332, 1485			-- fanout(506)
			, 31, 1504			-- fanout(507)
			, 755, 446			-- fanout(508)
			, 334			-- fanout(509)
			, 329, 1485			-- fanout(510)
			, 943, 480			-- fanout(511)
			, 313, 509			-- fanout(512)
			, 325, 1485			-- fanout(513)
			, 247, 1484			-- fanout(514)
			, 451			-- fanout(515)
			, 78			-- fanout(516)
			, 324, 1485			-- fanout(517)
			, 1171, 454			-- fanout(518)
			, 319, 481			-- fanout(519)
			, 321, 1485			-- fanout(520)
			, 1319, 541			-- fanout(521)
			, 547			-- fanout(522)
			, 1482, 531			-- fanout(523)
			, 340, 538			-- fanout(524)
			, 587, 545			-- fanout(525)
			, 1373, 837			-- fanout(526)
			, 177, 835			-- fanout(527)
			, 1409, 526			-- fanout(528)
			, 379, 842			-- fanout(529)
			, 548			-- fanout(530)
			, 1475, 827			-- fanout(531)
			, 350, 832			-- fanout(532)
			, 170, 838			-- fanout(533)
			, 164, 876			-- fanout(534)
			, 351, 799			-- fanout(535)
			, 347			-- fanout(536)
			, 630, 12			-- fanout(537)
			, 354			-- fanout(538)
			, 1383, 891			-- fanout(539)
			, 341, 536			-- fanout(540)
			, 166, 1240			-- fanout(541)
			, 336, 532			-- fanout(542)
			, 618, 12			-- fanout(543)
			, 337, 1228			-- fanout(544)
			, 594			-- fanout(545)
			, 338, 797			-- fanout(546)
			, 829			-- fanout(547)
			, 840			-- fanout(548)
			, 667, 38			-- fanout(549)
			, 1404, 853			-- fanout(550)
			, 1495, 843			-- fanout(551)
			, 668, 38			-- fanout(552)
			, 1406, 857			-- fanout(553)
			, 684, 38			-- fanout(554)
			, 847			-- fanout(555)
			, 1395, 851			-- fanout(556)
			, 1432, 863			-- fanout(557)
			, 1403, 855			-- fanout(558)
			, 1501, 551			-- fanout(559)
			, 1399, 866			-- fanout(560)
			, 28, 35			-- fanout(561)
			, 1414, 802			-- fanout(562)
			, 375, 213			-- fanout(563)
			, 1415, 816			-- fanout(564)
			, 1412, 826			-- fanout(565)
			, 1418, 820			-- fanout(566)
			, 383, 544			-- fanout(567)
			, 1408, 822			-- fanout(568)
			, 1391, 860			-- fanout(569)
			, 1393, 823			-- fanout(570)
			, 634, 1330			-- fanout(571)
			, 1413, 825			-- fanout(572)
			, 1392, 565			-- fanout(573)
			, 1424, 872			-- fanout(574)
			, 395, 881			-- fanout(575)
			, 1421, 885			-- fanout(576)
			, 1371, 874			-- fanout(577)
			, 20, 35			-- fanout(578)
			, 399, 1283			-- fanout(579)
			, 1475, 875			-- fanout(580)
			, 656, 38			-- fanout(581)
			, 1451, 576			-- fanout(582)
			, 1447, 871			-- fanout(583)
			, 426, 870			-- fanout(584)
			, 1450, 592			-- fanout(585)
			, 588			-- fanout(586)
			, 1472, 594			-- fanout(587)
			, 26			-- fanout(588)
			, 649, 38			-- fanout(589)
			, 555			-- fanout(590)
			, 659, 38			-- fanout(591)
			, 1420			-- fanout(592)
			, 673, 38			-- fanout(593)
			, 1464, 892			-- fanout(594)
			, 651, 849			-- fanout(595)
			, 652, 38			-- fanout(596)
			, 1407, 556			-- fanout(597)
			, 653, 38			-- fanout(598)
			, 422, 542			-- fanout(599)
			, 1436, 606			-- fanout(600)
			, 445, 599			-- fanout(601)
			, 1389, 605			-- fanout(602)
			, 522			-- fanout(603)
			, 1443, 86			-- fanout(604)
			, 1381, 534			-- fanout(605)
			, 1463, 539			-- fanout(606)
			, 1462, 889			-- fanout(607)
			, 1247, 1097			-- fanout(608)
			, 1456, 583			-- fanout(609)
			, 1445, 574			-- fanout(610)
			, 1482, 580			-- fanout(611)
			, 417, 579			-- fanout(612)
			, 1379, 577			-- fanout(613)
			, 1468, 573			-- fanout(614)
			, 1471, 683			-- fanout(615)
			, 438, 627			-- fanout(616)
			, 1494, 614			-- fanout(617)
			, 1417, 96			-- fanout(618)
			, 1430			-- fanout(619)
			, 376, 571			-- fanout(620)
			, 603			-- fanout(621)
			, 1170, 559			-- fanout(622)
			, 1407, 629			-- fanout(623)
			, 437, 535			-- fanout(624)
			, 1182			-- fanout(625)
			, 1403, 527			-- fanout(626)
			, 434, 567			-- fanout(627)
			, 1045, 61			-- fanout(628)
			, 1395, 521			-- fanout(629)
			, 1375, 96			-- fanout(630)
			, 1466, 86			-- fanout(631)
			, 204			-- fanout(632)
			, 467, 81			-- fanout(633)
			, 1043, 1458			-- fanout(634)
			, 586			-- fanout(635)
			, 1482, 640			-- fanout(636)
			, 487			-- fanout(637)
			, 1081, 628			-- fanout(638)
			, 359			-- fanout(639)
			, 1475, 597			-- fanout(640)
			, 366, 639			-- fanout(641)
			, 1485, 560			-- fanout(642)
			, 1502, 615			-- fanout(643)
			, 904			-- fanout(644)
			, 1008, 676			-- fanout(645)
			, 1133, 600			-- fanout(646)
			, 910, 1441			-- fanout(647)
			, 908, 760			-- fanout(648)
			, 1242, 122			-- fanout(649)
			, 914, 191			-- fanout(650)
			, 1309, 608			-- fanout(651)
			, 1204, 122			-- fanout(652)
			, 1246, 122			-- fanout(653)
			, 1464, 602			-- fanout(654)
			, 429, 660			-- fanout(655)
			, 1240, 122			-- fanout(656)
			, 1164, 646			-- fanout(657)
			, 913, 773			-- fanout(658)
			, 1236, 122			-- fanout(659)
			, 428			-- fanout(660)
			, 511, 672			-- fanout(661)
			, 922, 201			-- fanout(662)
			, 916, 1460			-- fanout(663)
			, 1459, 678			-- fanout(664)
			, 926, 790			-- fanout(665)
			, 490			-- fanout(666)
			, 1216, 122			-- fanout(667)
			, 1211, 122			-- fanout(668)
			, 1134, 582			-- fanout(669)
			, 489, 633			-- fanout(670)
			, 925, 1473			-- fanout(671)
			, 480, 612			-- fanout(672)
			, 1199, 122			-- fanout(673)
			, 1126, 130			-- fanout(674)
			, 928, 218			-- fanout(675)
			, 989, 102			-- fanout(676)
			, 476, 575			-- fanout(677)
			, 1442, 613			-- fanout(678)
			, 398, 595			-- fanout(679)
			, 1129, 669			-- fanout(680)
			, 478, 666			-- fanout(681)
			, 635			-- fanout(682)
			, 1142, 130			-- fanout(683)
			, 1206, 122			-- fanout(684)
			, 502, 176			-- fanout(685)
			, 1193, 689			-- fanout(686)
			, 455			-- fanout(687)
			, 1482, 696			-- fanout(688)
			, 1148			-- fanout(689)
			, 1190, 368			-- fanout(690)
			, 419, 695			-- fanout(691)
			, 198, 616			-- fanout(692)
			, 240			-- fanout(693)
			, 1158			-- fanout(694)
			, 411			-- fanout(695)
			, 1475, 623			-- fanout(696)
			, 514, 176			-- fanout(697)
			, 1155, 701			-- fanout(698)
			, 217			-- fanout(699)
			, 1472, 654			-- fanout(700)
			, 1166			-- fanout(701)
			, 1382, 1113			-- fanout(702)
			, 1407, 709			-- fanout(703)
			, 642, 1034			-- fanout(704)
			, 528, 714			-- fanout(705)
			, 1388, 1044			-- fanout(706)
			, 66, 1122			-- fanout(707)
			, 543, 498			-- fanout(708)
			, 1395, 1057			-- fanout(709)
			, 1397, 706			-- fanout(710)
			, 1274			-- fanout(711)
			, 79, 611			-- fanout(712)
			, 1403, 1067			-- fanout(713)
			, 526, 1056			-- fanout(714)
			, 74, 587			-- fanout(715)
			, 610			-- fanout(716)
			, 1082			-- fanout(717)
			, 47, 1073			-- fanout(718)
			, 48, 747			-- fanout(719)
			, 554, 213			-- fanout(720)
			, 1319, 740			-- fanout(721)
			, 1482, 736			-- fanout(722)
			, 552, 213			-- fanout(723)
			, 549, 213			-- fanout(724)
			, 598, 213			-- fanout(725)
			, 743			-- fanout(726)
			, 10, 1075			-- fanout(727)
			, 785, 1091			-- fanout(728)
			, 596, 213			-- fanout(729)
			, 91, 718			-- fanout(730)
			, 93, 748			-- fanout(731)
			, 50, 745			-- fanout(732)
			, 264, 1077			-- fanout(733)
			, 593, 213			-- fanout(734)
			, 177, 1092			-- fanout(735)
			, 1475, 1086			-- fanout(736)
			, 4			-- fanout(737)
			, 819, 1064			-- fanout(738)
			, 167, 1043			-- fanout(739)
			, 166, 1446			-- fanout(740)
			, 571, 0			-- fanout(741)
			, 1046			-- fanout(742)
			, 1443			-- fanout(743)
			, 296, 733			-- fanout(744)
			, 46			-- fanout(745)
			, 71			-- fanout(746)
			, 45, 1081			-- fanout(747)
			, 70, 1455			-- fanout(748)
			, 79, 636			-- fanout(749)
			, 140, 1496			-- fanout(750)
			, 1403, 1107			-- fanout(751)
			, 583, 1124			-- fanout(752)
			, 1395, 1099			-- fanout(753)
			, 81, 226			-- fanout(754)
			, 515, 1096			-- fanout(755)
			, 76, 1303			-- fanout(756)
			, 1442, 1104			-- fanout(757)
			, 114, 226			-- fanout(758)
			, 609, 752			-- fanout(759)
			, 188			-- fanout(760)
			, 610, 769			-- fanout(761)
			, 1437, 1103			-- fanout(762)
			, 595, 1070			-- fanout(763)
			, 591, 213			-- fanout(764)
			, 589, 213			-- fanout(765)
			, 95, 617			-- fanout(766)
			, 686			-- fanout(767)
			, 320, 1115			-- fanout(768)
			, 574, 1121			-- fanout(769)
			, 1466			-- fanout(770)
			, 581, 213			-- fanout(771)
			, 1441			-- fanout(772)
			, 333			-- fanout(773)
			, 1475, 703			-- fanout(774)
			, 103, 252			-- fanout(775)
			, 604, 245			-- fanout(776)
			, 1452, 702			-- fanout(777)
			, 711			-- fanout(778)
			, 177, 712			-- fanout(779)
			, 164, 750			-- fanout(780)
			, 545			-- fanout(781)
			, 348			-- fanout(782)
			, 108, 897			-- fanout(783)
			, 148, 707			-- fanout(784)
			, 169, 715			-- fanout(785)
			, 166, 1491			-- fanout(786)
			, 716			-- fanout(787)
			, 770			-- fanout(788)
			, 1460			-- fanout(789)
			, 156			-- fanout(790)
			, 1470, 710			-- fanout(791)
			, 101, 1490			-- fanout(792)
			, 1459, 757			-- fanout(793)
			, 1093, 1117			-- fanout(794)
			, 385			-- fanout(795)
			, 1407, 753			-- fanout(796)
			, 620, 741			-- fanout(797)
			, 1126			-- fanout(798)
			, 619, 50			-- fanout(799)
			, 1473			-- fanout(800)
			, 639			-- fanout(801)
			, 129, 746			-- fanout(802)
			, 726			-- fanout(803)
			, 172, 719			-- fanout(804)
			, 631, 245			-- fanout(805)
			, 1319, 786			-- fanout(806)
			, 1482, 774			-- fanout(807)
			, 142, 775			-- fanout(808)
			, 147, 792			-- fanout(809)
			, 1493, 471			-- fanout(810)
			, 18, 744			-- fanout(811)
			, 145, 657			-- fanout(812)
			, 525, 781			-- fanout(813)
			, 615, 856			-- fanout(814)
			, 166, 1197			-- fanout(815)
			, 162, 78			-- fanout(816)
			, 561, 281			-- fanout(817)
			, 161, 766			-- fanout(818)
			, 883, 728			-- fanout(819)
			, 163, 974			-- fanout(820)
			, 1416, 268			-- fanout(821)
			, 153			-- fanout(822)
			, 1338, 963			-- fanout(823)
			, 3			-- fanout(824)
			, 1341, 686			-- fanout(825)
			, 1337, 831			-- fanout(826)
			, 1407, 841			-- fanout(827)
			, 183, 804			-- fanout(828)
			, 798			-- fanout(829)
			, 641, 801			-- fanout(830)
			, 181, 1167			-- fanout(831)
			, 643, 814			-- fanout(832)
			, 742			-- fanout(833)
			, 178, 731			-- fanout(834)
			, 79, 688			-- fanout(835)
			, 1403, 735			-- fanout(836)
			, 152, 834			-- fanout(837)
			, 75, 72			-- fanout(838)
			, 186, 261			-- fanout(839)
			, 803			-- fanout(840)
			, 1395, 721			-- fanout(841)
			, 632, 344			-- fanout(842)
			, 1431, 821			-- fanout(843)
			, 655, 862			-- fanout(844)
			, 1328, 1217			-- fanout(845)
			, 124, 1206			-- fanout(846)
			, 858			-- fanout(847)
			, 1381, 780			-- fanout(848)
			, 608, 1006			-- fanout(849)
			, 701			-- fanout(850)
			, 1319, 815			-- fanout(851)
			, 1482, 864			-- fanout(852)
			, 1343, 996			-- fanout(853)
			, 674, 279			-- fanout(854)
			, 177, 749			-- fanout(855)
			, 683, 279			-- fanout(856)
			, 1346, 348			-- fanout(857)
			, 788			-- fanout(858)
			, 679, 763			-- fanout(859)
			, 1335, 106			-- fanout(860)
			, 168, 756			-- fanout(861)
			, 660			-- fanout(862)
			, 1321, 385			-- fanout(863)
			, 1475, 796			-- fanout(864)
			, 578, 281			-- fanout(865)
			, 1342, 149			-- fanout(866)
			, 1355, 888			-- fanout(867)
			, 687			-- fanout(868)
			, 1358, 812			-- fanout(869)
			, 693, 401			-- fanout(870)
			, 1356, 887			-- fanout(871)
			, 1348, 880			-- fanout(872)
			, 356, 868			-- fanout(873)
			, 139, 846			-- fanout(874)
			, 1407, 879			-- fanout(875)
			, 140, 1246			-- fanout(876)
			, 349, 886			-- fanout(877)
			, 778			-- fanout(878)
			, 1395, 806			-- fanout(879)
			, 1366, 809			-- fanout(880)
			, 699, 362			-- fanout(881)
			, 698, 850			-- fanout(882)
			, 1403, 779			-- fanout(883)
			, 695			-- fanout(884)
			, 1353, 845			-- fanout(885)
			, 694			-- fanout(886)
			, 1347, 808			-- fanout(887)
			, 1369			-- fanout(888)
			, 1370, 783			-- fanout(889)
			, 691, 884			-- fanout(890)
			, 1352, 1207			-- fanout(891)
			, 1389, 848			-- fanout(892)
			, 1051, 338			-- fanout(893)
			, 1334, 1233			-- fanout(894)
			, 234, 1305			-- fanout(895)
			, 67, 793			-- fanout(896)
			, 235, 920			-- fanout(897)
			, 231, 917			-- fanout(898)
			, 190, 911			-- fanout(899)
			, 1306			-- fanout(900)
			, 738, 1262			-- fanout(901)
			, 742, 1269			-- fanout(902)
			, 307			-- fanout(903)
			, 822			-- fanout(904)
			, 1319, 919			-- fanout(905)
			, 1065, 338			-- fanout(906)
			, 233, 918			-- fanout(907)
			, 820, 1435			-- fanout(908)
			, 1249			-- fanout(909)
			, 816, 516			-- fanout(910)
			, 508, 1268			-- fanout(911)
			, 716, 761			-- fanout(912)
			, 823, 1448			-- fanout(913)
			, 825, 767			-- fanout(914)
			, 177, 1227			-- fanout(915)
			, 860, 195			-- fanout(916)
			, 229, 1266			-- fanout(917)
			, 225, 1275			-- fanout(918)
			, 166, 94			-- fanout(919)
			, 242			-- fanout(920)
			, 241, 1232			-- fanout(921)
			, 857, 782			-- fanout(922)
			, 245, 1276			-- fanout(923)
			, 246			-- fanout(924)
			, 866, 207			-- fanout(925)
			, 853, 1467			-- fanout(926)
			, 1084, 935			-- fanout(927)
			, 863, 795			-- fanout(928)
			, 981, 1265			-- fanout(929)
			, 730, 950			-- fanout(930)
			, 731, 944			-- fanout(931)
			, 269			-- fanout(932)
			, 249, 1298			-- fanout(933)
			, 1407, 941			-- fanout(934)
			, 1048			-- fanout(935)
			, 267, 933			-- fanout(936)
			, 79, 807			-- fanout(937)
			, 1403, 1297			-- fanout(938)
			, 1091, 813			-- fanout(939)
			, 203, 1286			-- fanout(940)
			, 1395, 1288			-- fanout(941)
			, 200, 951			-- fanout(942)
			, 909			-- fanout(943)
			, 748, 114			-- fanout(944)
			, 669, 1287			-- fanout(945)
			, 254, 1252			-- fanout(946)
			, 244, 946			-- fanout(947)
			, 194, 123			-- fanout(948)
			, 717, 1259			-- fanout(949)
			, 718, 1299			-- fanout(950)
			, 193, 1250			-- fanout(951)
			, 1106			-- fanout(952)
			, 1482, 962			-- fanout(953)
			, 967			-- fanout(954)
			, 54, 398			-- fanout(955)
			, 680			-- fanout(956)
			, 292, 959			-- fanout(957)
			, 223, 1301			-- fanout(958)
			, 262			-- fanout(959)
			, 177, 1315			-- fanout(960)
			, 1118			-- fanout(961)
			, 1475, 1312			-- fanout(962)
			, 260, 966			-- fanout(963)
			, 1117, 1317			-- fanout(964)
			, 272, 932			-- fanout(965)
			, 257			-- fanout(966)
			, 1311			-- fanout(967)
			, 166, 134			-- fanout(968)
			, 206, 948			-- fanout(969)
			, 657			-- fanout(970)
			, 1080, 975			-- fanout(971)
			, 342, 1049			-- fanout(972)
			, 158, 1281			-- fanout(973)
			, 274, 924			-- fanout(974)
			, 1074			-- fanout(975)
			, 216, 940			-- fanout(976)
			, 255, 1037			-- fanout(977)
			, 280, 895			-- fanout(978)
			, 79, 852			-- fanout(979)
			, 1403, 915			-- fanout(980)
			, 279, 1304			-- fanout(981)
			, 781			-- fanout(982)
			, 787, 912			-- fanout(983)
			, 1395, 905			-- fanout(984)
			, 275, 1009			-- fanout(985)
			, 1281, 250			-- fanout(986)
			, 282, 898			-- fanout(987)
			, 900			-- fanout(988)
			, 112, 407			-- fanout(989)
			, 809, 994			-- fanout(990)
			, 189, 1052			-- fanout(991)
			, 808, 1003			-- fanout(992)
			, 124, 1345			-- fanout(993)
			, 792, 186			-- fanout(994)
			, 1434, 894			-- fanout(995)
			, 277, 1002			-- fanout(996)
			, 364, 972			-- fanout(997)
			, 94, 398			-- fanout(998)
			, 236, 626			-- fanout(999)
			, 291, 977			-- fanout(1000)
			, 65, 1143			-- fanout(1001)
			, 283			-- fanout(1002)
			, 775, 400			-- fanout(1003)
			, 568, 904			-- fanout(1004)
			, 1119, 952			-- fanout(1005)
			, 1097, 961			-- fanout(1006)
			, 1319, 968			-- fanout(1007)
			, 128, 989			-- fanout(1008)
			, 295			-- fanout(1009)
			, 778, 1307			-- fanout(1010)
			, 125, 416			-- fanout(1011)
			, 566, 908			-- fanout(1012)
			, 1042			-- fanout(1013)
			, 326, 1061			-- fanout(1014)
			, 572, 914			-- fanout(1015)
			, 564, 910			-- fanout(1016)
			, 1475, 934			-- fanout(1017)
			, 570, 913			-- fanout(1018)
			, 199, 991			-- fanout(1019)
			, 833, 902			-- fanout(1020)
			, 166, 1322			-- fanout(1021)
			, 327, 437			-- fanout(1022)
			, 834, 931			-- fanout(1023)
			, 302, 642			-- fanout(1024)
			, 569, 916			-- fanout(1025)
			, 550, 926			-- fanout(1026)
			, 553, 922			-- fanout(1027)
			, 560, 925			-- fanout(1028)
			, 988			-- fanout(1029)
			, 154, 1011			-- fanout(1030)
			, 144, 421			-- fanout(1031)
			, 813, 982			-- fanout(1032)
			, 157, 896			-- fanout(1033)
			, 557, 928			-- fanout(1034)
			, 304, 978			-- fanout(1035)
			, 306, 987			-- fanout(1036)
			, 298, 437			-- fanout(1037)
			, 1407, 984			-- fanout(1038)
			, 8, 1014			-- fanout(1039)
			, 1098			-- fanout(1040)
			, 139, 993			-- fanout(1041)
			, 943			-- fanout(1042)
			, 69, 284			-- fanout(1043)
			, 173, 1031			-- fanout(1044)
			, 315, 452			-- fanout(1045)
			, 867			-- fanout(1046)
			, 179, 471			-- fanout(1047)
			, 64			-- fanout(1048)
			, 171, 471			-- fanout(1049)
			, 184, 471			-- fanout(1050)
			, 1457, 442			-- fanout(1051)
			, 182, 471			-- fanout(1052)
			, 1324, 471			-- fanout(1053)
			, 331, 936			-- fanout(1054)
			, 1318, 471			-- fanout(1055)
			, 837, 1023			-- fanout(1056)
			, 1319, 1021			-- fanout(1057)
			, 1482, 1017			-- fanout(1058)
			, 220, 464			-- fanout(1059)
			, 261, 958			-- fanout(1060)
			, 1329, 471			-- fanout(1061)
			, 311, 1054			-- fanout(1062)
			, 817, 463			-- fanout(1063)
			, 728, 939			-- fanout(1064)
			, 1446, 442			-- fanout(1065)
			, 265, 969			-- fanout(1066)
			, 177, 937			-- fanout(1067)
			, 1327, 471			-- fanout(1068)
			, 160, 1001			-- fanout(1069)
			, 849, 1218			-- fanout(1070)
			, 1331, 471			-- fanout(1071)
			, 166, 1417			-- fanout(1072)
			, 5, 1083			-- fanout(1073)
			, 44			-- fanout(1074)
			, 289, 1066			-- fanout(1075)
			, 880, 990			-- fanout(1076)
			, 215, 1059			-- fanout(1077)
			, 878, 1010			-- fanout(1078)
			, 26, 476			-- fanout(1079)
			, 90, 1074			-- fanout(1080)
			, 13, 1045			-- fanout(1081)
			, 528			-- fanout(1082)
			, 14, 1000			-- fanout(1083)
			, 49, 1048			-- fanout(1084)
			, 865, 463			-- fanout(1085)
			, 1407, 1090			-- fanout(1086)
			, 17			-- fanout(1087)
			, 441, 997			-- fanout(1088)
			, 0, 1087			-- fanout(1089)
			, 1395, 1007			-- fanout(1090)
			, 715, 525			-- fanout(1091)
			, 79, 523			-- fanout(1092)
			, 1403, 960			-- fanout(1093)
			, 1112			-- fanout(1094)
			, 1359, 1008			-- fanout(1095)
			, 451, 1088			-- fanout(1096)
			, 1326, 1118			-- fanout(1097)
			, 19, 1110			-- fanout(1098)
			, 1319, 1072			-- fanout(1099)
			, 1482, 1114			-- fanout(1100)
			, 1138			-- fanout(1101)
			, 253, 1019			-- fanout(1102)
			, 1372, 1095			-- fanout(1103)
			, 1379, 1120			-- fanout(1104)
			, 537, 498			-- fanout(1105)
			, 84			-- fanout(1106)
			, 177, 979			-- fanout(1107)
			, 888			-- fanout(1108)
			, 887, 992			-- fanout(1109)
			, 30, 1035			-- fanout(1110)
			, 794, 964			-- fanout(1111)
			, 1029			-- fanout(1112)
			, 1376, 1030			-- fanout(1113)
			, 1475, 1038			-- fanout(1114)
			, 256, 1102			-- fanout(1115)
			, 25, 476			-- fanout(1116)
			, 973, 986			-- fanout(1117)
			, 1340			-- fanout(1118)
			, 72, 1106			-- fanout(1119)
			, 1371, 1041			-- fanout(1120)
			, 872, 1076			-- fanout(1121)
			, 53, 1039			-- fanout(1122)
			, 867, 1108			-- fanout(1123)
			, 871, 1109			-- fanout(1124)
			, 341			-- fanout(1125)
			, 906, 546			-- fanout(1126)
			, 99			-- fanout(1127)
			, 400, 562			-- fanout(1128)
			, 907, 1134			-- fanout(1129)
			, 396, 1139			-- fanout(1130)
			, 957			-- fanout(1131)
			, 985			-- fanout(1132)
			, 946, 1436			-- fanout(1133)
			, 918, 1451			-- fanout(1134)
			, 698			-- fanout(1135)
			, 1419			-- fanout(1136)
			, 80			-- fanout(1137)
			, 401, 1479			-- fanout(1138)
			, 377, 1157			-- fanout(1139)
			, 391, 1486			-- fanout(1140)
			, 349			-- fanout(1141)
			, 893, 546			-- fanout(1142)
			, 200, 1487			-- fanout(1143)
			, 79, 953			-- fanout(1144)
			, 119			-- fanout(1145)
			, 965			-- fanout(1146)
			, 939, 1032			-- fanout(1147)
			, 932			-- fanout(1148)
			, 358, 1165			-- fanout(1149)
			, 504, 1453			-- fanout(1150)
			, 1294, 1476			-- fanout(1151)
			, 1289			-- fanout(1152)
			, 1474			-- fanout(1153)
			, 52			-- fanout(1154)
			, 927, 1166			-- fanout(1155)
			, 360, 1199			-- fanout(1156)
			, 423, 558			-- fanout(1157)
			, 975			-- fanout(1158)
			, 420, 278			-- fanout(1159)
			, 448, 1163			-- fanout(1160)
			, 447, 151			-- fanout(1161)
			, 617			-- fanout(1162)
			, 430, 276			-- fanout(1163)
			, 947, 1133			-- fanout(1164)
			, 343, 1216			-- fanout(1165)
			, 935			-- fanout(1166)
			, 410, 562			-- fanout(1167)
			, 957, 1196			-- fanout(1168)
			, 952			-- fanout(1169)
			, 439, 1501			-- fanout(1170)
			, 987, 1481			-- fanout(1171)
			, 964, 1499			-- fanout(1172)
			, 440, 1062			-- fanout(1173)
			, 1502			-- fanout(1174)
			, 961			-- fanout(1175)
			, 1174			-- fanout(1176)
			, 79, 1058			-- fanout(1177)
			, 1009			-- fanout(1178)
			, 1232, 1040			-- fanout(1179)
			, 1000, 1190			-- fanout(1180)
			, 1380, 1478			-- fanout(1181)
			, 473, 1170			-- fanout(1182)
			, 1005, 1169			-- fanout(1183)
			, 374, 1156			-- fanout(1184)
			, 1036			-- fanout(1185)
			, 327			-- fanout(1186)
			, 845, 310			-- fanout(1187)
			, 1465			-- fanout(1188)
			, 971, 1158			-- fanout(1189)
			, 977, 1239			-- fanout(1190)
			, 377, 1242			-- fanout(1191)
			, 1300, 1152			-- fanout(1192)
			, 965, 1148			-- fanout(1193)
			, 861, 1469			-- fanout(1194)
			, 432, 1159			-- fanout(1195)
			, 959			-- fanout(1196)
			, 425, 558			-- fanout(1197)
			, 1146			-- fanout(1198)
			, 409, 626			-- fanout(1199)
			, 1186			-- fanout(1200)
			, 885, 1187			-- fanout(1201)
			, 466, 1130			-- fanout(1202)
			, 1497			-- fanout(1203)
			, 416, 626			-- fanout(1204)
			, 1135			-- fanout(1205)
			, 415, 626			-- fanout(1206)
			, 457, 607			-- fanout(1207)
			, 1137			-- fanout(1208)
			, 485, 1223			-- fanout(1209)
			, 1141			-- fanout(1210)
			, 407, 626			-- fanout(1211)
			, 713, 1492			-- fanout(1212)
			, 177, 1144			-- fanout(1213)
			, 1145			-- fanout(1214)
			, 869, 1503			-- fanout(1215)
			, 404, 626			-- fanout(1216)
			, 475, 607			-- fanout(1217)
			, 1006, 1175			-- fanout(1218)
			, 1062			-- fanout(1219)
			, 166, 330			-- fanout(1220)
			, 396, 1191			-- fanout(1221)
			, 1489			-- fanout(1222)
			, 461, 1140			-- fanout(1223)
			, 985, 1178			-- fanout(1224)
			, 481, 31			-- fanout(1225)
			, 510, 642			-- fanout(1226)
			, 79, 1100			-- fanout(1227)
			, 1022, 624			-- fanout(1228)
			, 506, 642			-- fanout(1229)
			, 509			-- fanout(1230)
			, 503, 1160			-- fanout(1231)
			, 483, 1098			-- fanout(1232)
			, 118, 1101			-- fanout(1233)
			, 226, 1150			-- fanout(1234)
			, 1125			-- fanout(1235)
			, 421, 626			-- fanout(1236)
			, 1127			-- fanout(1237)
			, 474, 1202			-- fanout(1238)
			, 1037, 624			-- fanout(1239)
			, 425, 626			-- fanout(1240)
			, 1131			-- fanout(1241)
			, 423, 626			-- fanout(1242)
			, 482, 449			-- fanout(1243)
			, 1319, 1220			-- fanout(1244)
			, 1132			-- fanout(1245)
			, 418, 626			-- fanout(1246)
			, 56, 1326			-- fanout(1247)
			, 1153			-- fanout(1248)
			, 1264			-- fanout(1249)
			, 460, 1253			-- fanout(1250)
			, 501, 1195			-- fanout(1251)
			, 196, 1251			-- fanout(1252)
			, 453, 1184			-- fanout(1253)
			, 491, 642			-- fanout(1254)
			, 166, 20			-- fanout(1255)
			, 499, 22			-- fanout(1256)
			, 500, 642			-- fanout(1257)
			, 1087			-- fanout(1258)
			, 1082, 705			-- fanout(1259)
			, 1083, 1180			-- fanout(1260)
			, 513, 642			-- fanout(1261)
			, 1064, 1147			-- fanout(1262)
			, 497, 642			-- fanout(1263)
			, 25			-- fanout(1264)
			, 921, 1179			-- fanout(1265)
			, 519, 1225			-- fanout(1266)
			, 492, 642			-- fanout(1267)
			, 446, 1272			-- fanout(1268)
			, 1046, 1123			-- fanout(1269)
			, 520, 642			-- fanout(1270)
			, 143, 1154			-- fanout(1271)
			, 435, 1149			-- fanout(1272)
			, 517, 642			-- fanout(1273)
			, 512, 1230			-- fanout(1274)
			, 494, 1231			-- fanout(1275)
			, 493, 1161			-- fanout(1276)
			, 1079, 677			-- fanout(1277)
			, 1440			-- fanout(1278)
			, 1200			-- fanout(1279)
			, 576, 1201			-- fanout(1280)
			, 63, 462			-- fanout(1281)
			, 1111, 1172			-- fanout(1282)
			, 1116, 677			-- fanout(1283)
			, 998, 679			-- fanout(1284)
			, 222, 1209			-- fanout(1285)
			, 474, 1293			-- fanout(1286)
			, 582, 1280			-- fanout(1287)
			, 1319, 1255			-- fanout(1288)
			, 757			-- fanout(1289)
			, 1089, 1258			-- fanout(1290)
			, 955, 679			-- fanout(1291)
			, 1176			-- fanout(1292)
			, 466, 1221			-- fanout(1293)
			, 558, 1194			-- fanout(1294)
			, 202, 1173			-- fanout(1295)
			, 1292			-- fanout(1296)
			, 177, 1177			-- fanout(1297)
			, 192, 1256			-- fanout(1298)
			, 1073, 1260			-- fanout(1299)
			, 793, 1289			-- fanout(1300)
			, 465, 737			-- fanout(1301)
			, 607, 1215			-- fanout(1302)
			, 216, 1310			-- fanout(1303)
			, 238, 1243			-- fanout(1304)
			, 239, 92			-- fanout(1305)
			, 697			-- fanout(1306)
			, 711, 1450			-- fanout(1307)
			, 1235			-- fanout(1308)
			, 155, 1247			-- fanout(1309)
			, 203, 1238			-- fanout(1310)
			, 1279			-- fanout(1311)
			, 1407, 1313			-- fanout(1312)
			, 1395, 1244			-- fanout(1313)
			, 224, 1285			-- fanout(1314)
			, 79, 722			-- fanout(1315)
			, 1403, 1213			-- fanout(1316)
			, 986, 478			-- fanout(1317)
			, 1261, 704			-- fanout(1318)
			, 402, 166			-- fanout(1319)
			, 586, 159			-- fanout(1320)
			, 1132, 1224			-- fanout(1321)
			, 425, 713			-- fanout(1322)
			, 575, 115			-- fanout(1323)
			, 1263, 704			-- fanout(1324)
			, 1426			-- fanout(1325)
			, 190, 1340			-- fanout(1326)
			, 1254, 704			-- fanout(1327)
			, 1163, 475			-- fanout(1328)
			, 1267, 704			-- fanout(1329)
			, 1458, 1325			-- fanout(1330)
			, 1257, 704			-- fanout(1331)
			, 678			-- fanout(1332)
			, 360, 1378			-- fanout(1333)
			, 584, 118			-- fanout(1334)
			, 1141, 877			-- fanout(1335)
			, 416, 713			-- fanout(1336)
			, 1140, 181			-- fanout(1337)
			, 1145, 260			-- fanout(1338)
			, 1433, 1192			-- fanout(1339)
			, 508, 117			-- fanout(1340)
			, 1146, 1193			-- fanout(1341)
			, 1125, 540			-- fanout(1342)
			, 1127, 277			-- fanout(1343)
			, 579, 433			-- fanout(1344)
			, 415, 713			-- fanout(1345)
			, 1131, 1168			-- fanout(1346)
			, 142			-- fanout(1347)
			, 1366			-- fanout(1348)
			, 700, 1365			-- fanout(1349)
			, 1173, 1219			-- fanout(1350)
			, 603, 138			-- fanout(1351)
			, 1159, 457			-- fanout(1352)
			, 1160, 1328			-- fanout(1353)
			, 621, 1351			-- fanout(1354)
			, 1192, 1369			-- fanout(1355)
			, 1347			-- fanout(1356)
			, 601, 1367			-- fanout(1357)
			, 1188, 145			-- fanout(1358)
			, 733, 128			-- fanout(1359)
			, 612, 1344			-- fanout(1360)
			, 374, 1333			-- fanout(1361)
			, 664, 1332			-- fanout(1362)
			, 1151, 109			-- fanout(1363)
			, 1444, 738			-- fanout(1364)
			, 654			-- fanout(1365)
			, 147			-- fanout(1366)
			, 599, 150			-- fanout(1367)
			, 1438, 738			-- fanout(1368)
			, 1152			-- fanout(1369)
			, 1153, 108			-- fanout(1370)
			, 444, 139			-- fanout(1371)
			, 744, 1359			-- fanout(1372)
			, 152			-- fanout(1373)
			, 1469, 313			-- fanout(1374)
			, 418, 751			-- fanout(1375)
			, 551, 154			-- fanout(1376)
			, 818, 137			-- fanout(1377)
			, 409, 751			-- fanout(1378)
			, 454, 1371			-- fanout(1379)
			, 624, 135			-- fanout(1380)
			, 458, 164			-- fanout(1381)
			, 559, 1376			-- fanout(1382)
			, 1195, 1352			-- fanout(1383)
			, 696			-- fanout(1384)
			, 627, 126			-- fanout(1385)
			, 1225, 507			-- fanout(1386)
			, 616, 1385			-- fanout(1387)
			, 345, 173			-- fanout(1388)
			, 468, 1381			-- fanout(1389)
			, 688, 1384			-- fanout(1390)
			, 1210, 1335			-- fanout(1391)
			, 1209, 1412			-- fanout(1392)
			, 1214, 1338			-- fanout(1393)
			, 1492, 1339			-- fanout(1394)
			, 472, 1319			-- fanout(1395)
						-- fanout(1396)
			, 352, 1388			-- fanout(1397)
			, 134, 794			-- fanout(1398)
			, 1235, 1342			-- fanout(1399)
			, 58, 1278			-- fanout(1400)
			, 666			-- fanout(1401)
			, 175			-- fanout(1402)
			, 471, 177			-- fanout(1403)
			, 1237, 1343			-- fanout(1404)
			, 635, 1320			-- fanout(1405)
			, 1241, 1346			-- fanout(1406)
			, 479, 1395			-- fanout(1407)
			, 1222, 153			-- fanout(1408)
			, 1373			-- fanout(1409)
			, 1266, 1386			-- fanout(1410)
			, 141, 794			-- fanout(1411)
			, 1223, 1337			-- fanout(1412)
			, 1198, 1341			-- fanout(1413)
			, 1203, 129			-- fanout(1414)
			, 1205, 162			-- fanout(1415)
			, 633, 754			-- fanout(1416)
			, 425, 751			-- fanout(1417)
			, 1208, 163			-- fanout(1418)
			, 1314			-- fanout(1419)
			, 1230			-- fanout(1420)
			, 1231, 1353			-- fanout(1421)
			, 661, 1427			-- fanout(1422)
			, 460, 1428			-- fanout(1423)
			, 1348			-- fanout(1424)
			, 1295, 1350			-- fanout(1425)
			, 297			-- fanout(1426)
			, 672, 1360			-- fanout(1427)
			, 453, 1361			-- fanout(1428)
			, 682, 1405			-- fanout(1429)
			, 681, 1401			-- fanout(1430)
			, 670, 1416			-- fanout(1431)
			, 1245, 1321			-- fanout(1432)
			, 896, 1300			-- fanout(1433)
			, 677, 1323			-- fanout(1434)
			, 974			-- fanout(1435)
			, 1252, 1463			-- fanout(1436)
			, 811, 1372			-- fanout(1437)
			, 1488, 819			-- fanout(1438)
			, 692, 1387			-- fanout(1439)
			, 344, 1439			-- fanout(1440)
			, 824			-- fanout(1441)
			, 518, 1379			-- fanout(1442)
			, 1291, 859			-- fanout(1443)
			, 1491, 819			-- fanout(1444)
			, 1424			-- fanout(1445)
			, 425, 836			-- fanout(1446)
			, 1356			-- fanout(1447)
			, 963			-- fanout(1448)
			, 697, 833			-- fanout(1449)
			, 1274, 1420			-- fanout(1450)
			, 1275, 1421			-- fanout(1451)
			, 622, 1382			-- fanout(1452)
			, 413, 903			-- fanout(1453)
			, 562, 1377			-- fanout(1454)
			, 685, 833			-- fanout(1455)
			, 1447			-- fanout(1456)
			, 423, 836			-- fanout(1457)
			, 284, 1426			-- fanout(1458)
			, 191			-- fanout(1459)
			, 625			-- fanout(1460)
			, 416, 836			-- fanout(1461)
			, 1248, 1370			-- fanout(1462)
			, 1251, 1383			-- fanout(1463)
			, 197, 1389			-- fanout(1464)
			, 947			-- fanout(1465)
			, 1284, 859			-- fanout(1466)
			, 996			-- fanout(1467)
			, 1285, 1392			-- fanout(1468)
			, 756, 89			-- fanout(1469)
			, 431, 1397			-- fanout(1470)
			, 1142			-- fanout(1471)
			, 201			-- fanout(1472)
			, 443			-- fanout(1473)
			, 60			-- fanout(1474)
			, 208, 1407			-- fanout(1475)
			, 1194, 1374			-- fanout(1476)
			, 917, 1410			-- fanout(1477)
			, 120, 1400			-- fanout(1478)
			, 365, 1422			-- fanout(1479)
						-- fanout(1480)
			, 898, 1477			-- fanout(1481)
			, 218			-- fanout(1482)
			, 370, 1505			-- fanout(1483)
			, 1212, 1394			-- fanout(1484)
			, 1308, 1399			-- fanout(1485)
			, 367, 248			-- fanout(1486)
			, 193, 1423			-- fanout(1487)
			, 421, 883			-- fanout(1488)
						-- fanout(1489)
			, 357, 878			-- fanout(1490)
			, 425, 883			-- fanout(1491)
			, 1033, 1433			-- fanout(1492)
			, 1024, 704			-- fanout(1493)
			, 1314, 1468			-- fanout(1494)
			, 382, 1431			-- fanout(1495)
			, 418, 883			-- fanout(1496)
			, 1396			-- fanout(1497)
			, 388			-- fanout(1498)
			, 1317, 681			-- fanout(1499)
			, 362, 1498			-- fanout(1500)
			, 363, 1495			-- fanout(1501)
			, 1471			-- fanout(1502)
			, 812, 970			-- fanout(1503)
			, 923, 1425			-- fanout(1504)
			, 386, 1429			-- fanout(1505)
		),
		fanout_base => (0, 2, 3, 5, 7, 9, 10, 12, 14, 16, 18, 20, 22, 24, 26, 27, 29, 31, 32, 34, 36, 38, 40, 42, 44, 46, 48, 50, 52, 54, 56, 58, 60, 61, 62, 64, 66, 68, 70, 72, 74, 76, 78, 79, 80, 82, 84, 85, 86, 88, 90, 92, 94, 95, 97, 99, 101, 103, 105, 107, 109, 111, 113, 115, 117, 119, 121, 123, 125, 127, 129, 130, 131, 133, 134, 136, 138, 140, 142, 144, 146, 148, 150, 151, 152, 154, 156, 157, 159, 160, 162, 164, 165, 167, 168, 170, 172, 174, 175, 177, 179, 180, 181, 183, 184, 186, 188, 190, 191, 193, 195, 196, 198, 200, 201, 203, 205, 206, 208, 210, 212, 214, 216, 218, 220, 222, 224, 226, 228, 230, 232, 233, 235, 237, 238, 240, 242, 244, 246, 248, 250, 252, 254, 255, 257, 259, 261, 263, 264, 266, 268, 270, 272, 273, 274, 276, 278, 279, 281, 283, 285, 287, 289, 291, 293, 295, 297, 299, 301, 303, 305, 307, 309, 311, 313, 315, 316, 318, 320, 321, 323, 325, 327, 329, 331, 333, 335, 337, 339, 339, 341, 342, 343, 345, 347, 349, 350, 351, 353, 355, 357, 358, 359, 361, 363, 365, 367, 369, 370, 372, 374, 376, 377, 379, 381, 383, 385, 386, 388, 389, 391, 393, 395, 396, 398, 399, 400, 402, 404, 406, 408, 409, 411, 413, 414, 416, 418, 420, 422, 424, 426, 428, 430, 431, 432, 433, 435, 436, 438, 440, 442, 444, 446, 448, 450, 451, 452, 454, 455, 457, 459, 461, 463, 464, 465, 467, 469, 471, 473, 475, 476, 478, 479, 481, 483, 485, 487, 489, 491, 493, 495, 497, 499, 501, 502, 504, 506, 507, 509, 511, 513, 515, 516, 518, 520, 522, 523, 525, 527, 529, 531, 533, 534, 536, 538, 540, 542, 544, 546, 548, 550, 552, 554, 556, 558, 560, 562, 564, 566, 568, 570, 572, 574, 575, 577, 579, 581, 583, 585, 586, 588, 590, 592, 594, 595, 596, 597, 599, 601, 603, 605, 607, 609, 610, 612, 614, 616, 618, 619, 621, 623, 625, 626, 628, 629, 630, 632, 634, 636, 638, 639, 641, 643, 645, 647, 648, 650, 652, 653, 655, 657, 658, 660, 662, 664, 666, 668, 670, 672, 674, 675, 677, 679, 681, 683, 685, 687, 688, 690, 691, 693, 695, 696, 698, 700, 702, 703, 705, 707, 709, 711, 713, 715, 717, 719, 721, 723, 725, 727, 728, 730, 732, 733, 734, 736, 738, 740, 742, 744, 746, 748, 749, 751, 753, 755, 757, 759, 760, 762, 763, 765, 766, 768, 769, 771, 773, 775, 777, 778, 780, 782, 784, 785, 787, 788, 790, 792, 794, 796, 797, 799, 801, 802, 804, 806, 808, 809, 811, 813, 815, 817, 819, 820, 822, 824, 826, 828, 830, 832, 834, 836, 838, 840, 842, 844, 846, 848, 849, 851, 853, 855, 857, 859, 861, 863, 865, 866, 868, 869, 871, 873, 874, 876, 878, 880, 881, 883, 885, 887, 889, 891, 893, 894, 896, 897, 899, 901, 903, 905, 907, 908, 910, 912, 914, 916, 918, 919, 920, 922, 924, 926, 928, 930, 931, 933, 935, 937, 939, 941, 943, 945, 946, 948, 950, 952, 954, 956, 957, 959, 960, 962, 964, 966, 968, 970, 972, 973, 975, 976, 977, 979, 981, 983, 985, 987, 989, 990, 992, 994, 996, 998, 1000, 1002, 1004, 1006, 1008, 1010, 1012, 1014, 1016, 1018, 1020, 1022, 1024, 1026, 1028, 1030, 1032, 1034, 1036, 1038, 1040, 1042, 1044, 1046, 1048, 1050, 1051, 1053, 1054, 1056, 1057, 1059, 1060, 1062, 1064, 1066, 1068, 1070, 1072, 1074, 1076, 1078, 1080, 1081, 1083, 1085, 1087, 1089, 1091, 1093, 1095, 1097, 1099, 1101, 1103, 1105, 1107, 1109, 1111, 1112, 1114, 1115, 1117, 1119, 1121, 1122, 1124, 1126, 1128, 1130, 1132, 1134, 1135, 1137, 1139, 1140, 1142, 1143, 1145, 1146, 1148, 1150, 1152, 1154, 1155, 1157, 1159, 1161, 1163, 1165, 1167, 1169, 1171, 1173, 1175, 1177, 1179, 1181, 1183, 1185, 1186, 1188, 1190, 1192, 1194, 1196, 1197, 1199, 1201, 1203, 1205, 1207, 1209, 1211, 1213, 1215, 1217, 1219, 1221, 1223, 1225, 1227, 1228, 1230, 1232, 1234, 1236, 1237, 1239, 1240, 1242, 1244, 1246, 1247, 1248, 1249, 1251, 1253, 1255, 1256, 1258, 1259, 1261, 1263, 1265, 1267, 1269, 1271, 1273, 1275, 1277, 1278, 1280, 1282, 1284, 1286, 1287, 1288, 1290, 1292, 1294, 1296, 1298, 1300, 1302, 1304, 1305, 1307, 1309, 1311, 1313, 1315, 1317, 1319, 1321, 1323, 1325, 1326, 1328, 1330, 1332, 1334, 1335, 1336, 1338, 1339, 1340, 1342, 1344, 1346, 1348, 1350, 1352, 1354, 1356, 1358, 1360, 1362, 1364, 1366, 1367, 1369, 1371, 1373, 1375, 1377, 1379, 1380, 1382, 1384, 1385, 1387, 1388, 1389, 1391, 1393, 1395, 1397, 1398, 1400, 1402, 1403, 1404, 1406, 1408, 1410, 1412, 1413, 1414, 1415, 1416, 1418, 1420, 1422, 1424, 1425, 1427, 1429, 1430, 1432, 1433, 1434, 1436, 1437, 1439, 1441, 1443, 1445, 1447, 1449, 1451, 1453, 1455, 1457, 1459, 1461, 1463, 1465, 1467, 1469, 1471, 1473, 1474, 1476, 1477, 1479, 1481, 1483, 1485, 1486, 1488, 1490, 1492, 1493, 1495, 1497, 1499, 1501, 1503, 1505, 1506, 1508, 1510, 1512, 1514, 1516, 1518, 1519, 1521, 1523, 1524, 1526, 1528, 1530, 1532, 1534, 1536, 1538, 1539, 1541, 1543, 1545, 1546, 1548, 1550, 1552, 1554, 1556, 1557, 1559, 1561, 1563, 1565, 1567, 1569, 1571, 1573, 1575, 1576, 1578, 1580, 1582, 1584, 1586, 1587, 1589, 1590, 1592, 1593, 1595, 1597, 1599, 1601, 1603, 1605, 1607, 1609, 1611, 1613, 1615, 1616, 1618, 1620, 1621, 1622, 1624, 1626, 1628, 1630, 1631, 1633, 1635, 1637, 1639, 1641, 1643, 1645, 1647, 1649, 1651, 1652, 1654, 1656, 1658, 1659, 1661, 1663, 1665, 1667, 1669, 1671, 1673, 1674, 1676, 1678, 1679, 1681, 1683, 1685, 1687, 1689, 1691, 1693, 1694, 1696, 1698, 1700, 1702, 1704, 1706, 1708, 1710, 1711, 1713, 1714, 1716, 1717, 1719, 1721, 1722, 1724, 1725, 1727, 1729, 1731, 1733, 1734, 1735, 1737, 1739, 1740, 1742, 1744, 1746, 1748, 1749, 1751, 1753, 1755, 1757, 1759, 1761, 1762, 1764, 1766, 1768, 1770, 1772, 1773, 1775, 1777, 1779, 1781, 1783, 1785, 1787, 1789, 1791, 1793, 1795, 1797, 1799, 1800, 1802, 1804, 1806, 1808, 1810, 1812, 1813, 1815, 1817, 1819, 1820, 1822, 1824, 1826, 1828, 1830, 1832, 1834, 1836, 1838, 1840, 1842, 1844, 1846, 1848, 1850, 1851, 1853, 1855, 1857, 1859, 1861, 1863, 1865, 1867, 1869, 1871, 1872, 1874, 1875, 1877, 1879, 1881, 1882, 1884, 1885, 1887, 1889, 1891, 1893, 1895, 1897, 1899, 1901, 1903, 1905, 1907, 1909, 1911, 1913, 1915, 1917, 1919, 1921, 1923, 1925, 1927, 1929, 1931, 1933, 1935, 1936, 1938, 1940, 1942, 1944, 1946, 1948, 1950, 1951, 1953, 1955, 1957, 1959, 1960, 1962, 1964, 1966, 1968, 1970, 1972, 1973, 1975, 1977, 1979, 1981, 1983, 1985, 1986, 1988, 1990, 1992, 1994, 1995, 1997, 1998, 2000, 2002, 2004, 2005, 2007, 2009, 2011, 2013, 2015, 2016, 2018, 2020, 2022, 2024, 2026, 2028, 2029, 2031, 2032, 2034, 2036, 2038, 2039, 2040, 2042, 2044, 2045, 2046, 2047, 2049, 2051, 2053, 2054, 2056, 2058, 2060, 2061, 2062, 2064, 2065, 2067, 2069, 2071, 2072, 2073, 2074, 2076, 2078, 2080, 2081, 2083, 2085, 2087, 2088, 2090, 2092, 2094, 2095, 2097, 2099, 2100, 2102, 2104, 2106, 2108, 2109, 2110, 2111, 2113, 2114, 2116, 2118, 2120, 2122, 2124, 2126, 2127, 2128, 2130, 2131, 2133, 2135, 2137, 2139, 2141, 2143, 2145, 2146, 2148, 2149, 2151, 2152, 2154, 2156, 2157, 2159, 2160, 2162, 2164, 2165, 2167, 2168, 2170, 2172, 2174, 2175, 2177, 2179, 2181, 2183, 2184, 2186, 2188, 2189, 2191, 2193, 2195, 2197, 2199, 2201, 2203, 2204, 2206, 2208, 2210, 2212, 2213, 2215, 2216, 2218, 2220, 2222, 2223, 2225, 2227, 2229, 2230, 2232, 2234, 2235, 2236, 2238, 2240, 2242, 2244, 2246, 2248, 2250, 2252, 2253, 2255, 2257, 2259, 2261, 2263, 2264, 2266, 2268, 2270, 2272, 2274, 2276, 2278, 2280, 2282, 2284, 2286, 2288, 2290, 2291, 2292, 2294, 2296, 2298, 2300, 2302, 2304, 2306, 2308, 2310, 2311, 2313, 2315, 2316, 2318, 2320, 2322, 2323, 2325, 2327, 2329, 2331, 2333, 2335, 2337, 2339, 2341, 2342, 2344, 2345, 2347, 2349, 2350, 2352, 2354, 2356, 2358, 2360, 2362, 2364, 2366, 2368, 2370, 2372, 2374, 2376, 2377, 2379, 2381, 2383, 2385, 2387, 2389, 2390, 2392, 2394, 2396, 2398, 2400, 2402, 2404, 2406, 2408, 2410, 2412, 2414, 2416, 2418, 2419, 2420, 2422, 2424, 2426, 2428, 2430, 2432, 2434, 2435, 2437, 2439, 2441, 2443, 2445, 2447, 2449, 2451, 2452, 2453, 2455, 2457, 2458, 2460, 2462, 2464, 2465, 2467, 2469, 2471, 2473, 2475, 2477, 2479, 2481, 2483, 2485, 2486, 2488, 2490, 2492, 2494, 2496, 2498, 2500, 2502, 2504, 2506, 2508, 2508, 2510, 2512, 2514, 2516, 2517, 2518, 2520, 2522, 2524, 2526, 2528, 2530, 2531, 2533, 2535, 2537, 2539, 2541, 2543, 2545, 2547, 2549, 2550, 2551, 2553, 2555, 2557, 2558, 2560, 2561, 2563, 2565, 2567, 2569, 2571, 2573, 2575, 2577, 2578, 2580, 2582, 2584, 2586, 2588, 2589, 2591, 2593, 2595, 2596, 2598, 2599, 2600, 2602, 2604, 2606, 2608, 2610, 2612, 2614, 2615, 2617, 2619, 2620, 2621, 2623, 2625, 2627, 2629, 2630, 2632, 2633, 2635, 2637, 2639, 2640, 2641, 2642, 2643, 2645, 2647, 2649, 2651, 2653, 2653, 2655, 2656, 2658, 2660, 2662, 2664, 2666, 2668, 2668, 2670, 2672, 2674, 2676, 2678, 2680, 2682, 2683, 2684, 2686, 2688, 2690, 2691, 2693, 2695, ab_params.nb_transitions)
);
end package;